
module tests();
    
    supply0 gnd;
    supply1 vdd;



    initial begin
        
    end
endmodule


