
module calculator(input vdd, inout gnd);



endmodule


